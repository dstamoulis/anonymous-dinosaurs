library verilog;
use verilog.vl_types.all;
entity testbenchPPR is
end testbenchPPR;
