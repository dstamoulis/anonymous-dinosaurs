library verilog;
use verilog.vl_types.all;
entity testbenchFTCfunct is
end testbenchFTCfunct;
