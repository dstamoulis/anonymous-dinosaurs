library verilog;
use verilog.vl_types.all;
entity \muddlib07__fulladder\ is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        cout            : out    vl_logic;
        s               : out    vl_logic
    );
end \muddlib07__fulladder\;
