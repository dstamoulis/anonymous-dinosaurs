library verilog;
use verilog.vl_types.all;
entity testbenchCHECK is
end testbenchCHECK;
