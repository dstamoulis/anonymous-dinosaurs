library verilog;
use verilog.vl_types.all;
entity testbenchCPA is
end testbenchCPA;
