library verilog;
use verilog.vl_types.all;
entity \muddlib07__a2o1_1x\ is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        y               : out    vl_logic
    );
end \muddlib07__a2o1_1x\;
