library verilog;
use verilog.vl_types.all;
entity testbenchXNOR is
end testbenchXNOR;
