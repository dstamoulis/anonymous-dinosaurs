library verilog;
use verilog.vl_types.all;
entity testbenchFTC is
end testbenchFTC;
