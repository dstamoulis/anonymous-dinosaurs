library verilog;
use verilog.vl_types.all;
entity testbenchPPRfunct is
end testbenchPPRfunct;
