library verilog;
use verilog.vl_types.all;
entity testbenchCPAfunct is
end testbenchCPAfunct;
